tb.poke(.addr(`HELLO_WORLD_REG_ADDR), .data(32'b00110000000000000000000000000001), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
tb.poke(.addr(`HELLO_WORLD_REG_ADDR), .data(32'b00110000000000000000000000000001), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
tb.poke(.addr(`HELLO_WORLD_REG_ADDR), .data(32'b00110000000000000000000000000010), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
tb.poke(.addr(`HELLO_WORLD_REG_ADDR), .data(32'b00110000000000000000000000000011), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
tb.peek(.addr(`HELLO_WORLD_REG_ADDR), .data(rdata), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
if (rdata == 32'he0000000) $display ("TEST PASSED"); else $error ("TEST FAILED");
tb.poke(.addr(`HELLO_WORLD_REG_ADDR), .data(32'b01000000000000000000000000000001), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
tb.peek(.addr(`HELLO_WORLD_REG_ADDR), .data(rdata), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
if (rdata == 32'b01000000000000000000000000000001) $display ("TEST PASSED"); else $error ("TEST FAILED");
tb.poke(.addr(`HELLO_WORLD_REG_ADDR), .data(32'b01000000000000000000000000000010), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
tb.peek(.addr(`HELLO_WORLD_REG_ADDR), .data(rdata), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
if (rdata == 32'b01000000000000000000000000000010) $display ("TEST PASSED"); else $error ("TEST FAILED");
tb.peek(.addr(`HELLO_WORLD_REG_ADDR), .data(rdata), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
if (rdata == 32'b01110000000000000000000000000001) $display ("TEST PASSED"); else $error ("TEST FAILED");
tb.poke(.addr(`HELLO_WORLD_REG_ADDR), .data(32'b01000000000000000000000000000011), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
tb.peek(.addr(`HELLO_WORLD_REG_ADDR), .data(rdata), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
if (rdata == 32'b01000000000000000000000000000011) $display ("TEST PASSED"); else $error ("TEST FAILED");
tb.peek(.addr(`HELLO_WORLD_REG_ADDR), .data(rdata), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
if (rdata == 32'b01100000000000000000000000000001) $display ("TEST PASSED"); else $error ("TEST FAILED");
tb.peek(.addr(`HELLO_WORLD_REG_ADDR), .data(rdata), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));
if (rdata == 32'he0000000) $display ("TEST PASSED"); else $error ("TEST FAILED");
